module ex7;
  int arr[3] = '{1, 2, 3};
  initial $display("arr = %p", arr);
endmodule

output : arr = '{1, 2, 3}
