module power;
  initial begin
    $display("2**3 = %0d", 2**3);
  end
endmodule

output : 
# KERNEL: 2**3 = 8
# KERNEL: Simulation has finished.
