module m7;
  int i = 0;
  initial begin
    do begin
      $display("i = %0d", i);
      i--;
      
    end while (i < 3);
   
  end
  
endmodule

output :

# KERNEL: i = 0
# KERNEL: i = -1
# KERNEL: i = -2
# KERNEL: i = -3
# KERNEL: i = -4
# KERNEL: i = -5
# KERNEL: i = -6
# KERNEL: i = -7
# KERNEL: i = -8
# KERNEL: i = -9
# KERNEL: i = -10
# KERNEL: i = -11
# KERNEL: i = -12
# KERNEL: i = -13
# KERNEL: i = -14
# KERNEL: i = -15
# KERNEL: i = -16
# KERNEL: i = -17
# KERNEL: i = -18
# KERNEL: i = -19
# KERNEL: i = -20
# KERNEL: i = -21
# KERNEL: i = -22
# KERNEL: i = -23
# KERNEL: i = -24
# KERNEL: i = -25
# KERNEL: i = -26
# KERNEL: i = -27
# KERNEL: i = -28
# KERNEL: i = -29
# KERNEL: i = -30
# KERNEL: i = -31
# KERNEL: i = -32
# KERNEL: i = -33
# KERNEL: i = -34
# KERNEL: i = -35
# KERNEL: i = -36
# KERNEL: i = -37
# KERNEL: i = -38
# KERNEL: i = -39
# KERNEL: i = -40
# KERNEL: i = -41
# KERNEL: i = -42
# KERNEL: i = -43
# KERNEL: i = -44
# KERNEL: i = -45
# KERNEL: i = -46
# KERNEL: i = -47
# KERNEL: i = -48
# KERNEL: i = -49
# KERNEL: i = -50
# KERNEL: i = -51
# KERNEL: i = -52
# KERNEL: i = -53
# KERNEL: i = -54
# KERNEL: i = -55
# KERNEL: i = -56
# KERNEL: i = -57
# KERNEL: i = -58
# KERNEL: i = -59
# KERNEL: i = -60
# KERNEL: i = -61
# KERNEL: i = -62
# KERNEL: i = -63
# KERNEL: i = -64
# KERNEL: i = -65
# KERNEL: i = -66
# KERNEL: i = -67
# KERNEL: i = -68
# KERNEL: i = -69
# KERNEL: i = -70
# KERNEL: i = -71
# KERNEL: i = -72
# KERNEL: i = -73
# KERNEL: i = -74
# KERNEL: i = -75
# KERNEL: i = -76
# KERNEL: i = -77
# KERNEL: i = -78
# KERNEL: i = -79
# KERNEL: i = -80
# KERNEL: i = -81
# KERNEL: i = -82
# KERNEL: i = -83
# KERNEL: i = -84
# KERNEL: i = -85
# KERNEL: i = -86
# KERNEL: i = -87
# KERNEL: i = -88
# KERNEL: i = -89
# KERNEL: i = -90
# KERNEL: i = -91
# KERNEL: i = -92
# KERNEL: i = -93
# KERNEL: i = -94
# KERNEL: i = -95
# KERNEL: i = -96
# KERNEL: i = -97
# KERNEL: i = -98
# KERNEL: i = -99
# KERNEL: i = -100
# KERNEL: i = -101
# KERNEL: i = -102
# KERNEL: i = -103
# KERNEL: i = -104
# KERNEL: i = -105
# KERNEL: i = -106
# KERNEL: i = -107
# KERNEL: i = -108
# KERNEL: i = -109
# KERNEL: i = -110
# KERNEL: i = -111
# KERNEL: i = -112
# KERNEL: i = -113
# KERNEL: i = -114
# KERNEL: i = -115
# KERNEL: i = -116
# KERNEL: i = -117
# KERNEL: i = -118
# KERNEL: i = -119
# KERNEL: i = -120
# KERNEL: i = -121
# KERNEL: i = -122
# KERNEL: i = -123
# KERNEL: i = -124
# KERNEL: i = -125
# KERNEL: i = -126
# KERNEL: i = -127
# KERNEL: i = -128
# KERNEL: i = -129
# KERNEL: i = -130
# KERNEL: i = -131
# KERNEL: i = -132
# KERNEL: i = -133
# KERNEL: i = -134
# KERNEL: i = -135
# KERNEL: i = -136
# KERNEL: i = -137
# KERNEL: i = -138
# KERNEL: i = -139
# KERNEL: i = -140
# KERNEL: i = -141
# KERNEL: i = -142
# KERNEL: i = -143
# KERNEL: i = -144
# KERNEL: i = -145
# KERNEL: i = -146
# KERNEL: i = -147
# KERNEL: i = -148
# KERNEL: i = -149
# KERNEL: i = -150
# KERNEL: i = -151
# KERNEL: i = -152
# KERNEL: i = -153
# KERNEL: i = -154
# KERNEL: i = -155
# KERNEL: i = -156
# KERNEL: i = -157
# KERNEL: i = -158
# KERNEL: i = -159
# KERNEL: i = -160
# KERNEL: i = -161
# KERNEL: i = -162
# KERNEL: i = -163
# KERNEL: i = -164
# KERNEL: i = -165
# KERNEL: i = -166
# KERNEL: i = -167
# KERNEL: i = -168
# KERNEL: i = -169
# KERNEL: i = -170
# KERNEL: i = -171
# KERNEL: i = -172
# KERNEL: i = -173
# KERNEL: i = -174
# KERNEL: i = -175
# KERNEL: i = -176
# KERNEL: i = -177
# KERNEL: i = -178
# KERNEL: i = -179
# KERNEL: i = -180
# KERNEL: i = -181
# KERNEL: i = -182
# KERNEL: i = -183
# KERNEL: i = -184
# KERNEL: i = -185
# KERNEL: i = -186
# KERNEL: i = -187
# KERNEL: i = -188
# KERNEL: i = -189
# KERNEL: i = -190
# KERNEL: i = -191
# KERNEL: i = -192
# KERNEL: i = -193
# KERNEL: i = -194
# KERNEL: i = -195
# KERNEL: i = -196
# KERNEL: i = -197
# KERNEL: i = -198
# KERNEL: i = -199
# KERNEL: i = -200
# KERNEL: i = -201
# KERNEL: i = -202
# KERNEL: i = -203
# KERNEL: i = -204
# KERNEL: i = -205
# KERNEL: i = -206
# KERNEL: i = -207
# KERNEL: i = -208
# KERNEL: i = -209
# KERNEL: i = -210
# KERNEL: i = -211
# KERNEL: i = -212
# KERNEL: i = -213
# KERNEL: i = -214
# KERNEL: i = -215
# KERNEL: i = -216
# KERNEL: i = -217
# KERNEL: i = -218
# KERNEL: i = -219
# KERNEL: i = -220
# KERNEL: i = -221
# KERNEL: i = -222
# KERNEL: i = -223
# KERNEL: i = -224
# KERNEL: i = -225
# KERNEL: i = -226
# KERNEL: i = -227
# KERNEL: i = -228
# KERNEL: i = -229
# KERNEL: i = -230
# KERNEL: i = -231
# KERNEL: i = -232
# KERNEL: i = -233
# KERNEL: i = -234
# KERNEL: i = -235
# KERNEL: i = -236
# KERNEL: i = -237
# KERNEL: i = -238
# KERNEL: i = -239
# KERNEL: i = -240
# KERNEL: i = -241
# KERNEL: i = -242
# KERNEL: i = -243
# KERNEL: i = -244
# KERNEL: i = -245
# KERNEL: i = -246
# KERNEL: i = -247
# KERNEL: i = -248
# KERNEL: i = -249
# KERNEL: i = -250
# KERNEL: i = -251
# KERNEL: i = -252
# KERNEL: i = -253
# KERNEL: i = -254
# KERNEL: i = -255
# KERNEL: i = -256
# KERNEL: i = -257
# KERNEL: i = -258
# KERNEL: i = -259
# KERNEL: i = -260
# KERNEL: i = -261
# KERNEL: i = -262
# KERNEL: i = -263
# KERNEL: i = -264
# KERNEL: i = -265
# KERNEL: i = -266
# KERNEL: i = -267
# KERNEL: i = -268
# KERNEL: i = -269
# KERNEL: i = -270
# KERNEL: i = -271
# KERNEL: i = -272
# KERNEL: i = -273
# KERNEL: i = -274
# KERNEL: i = -275
# KERNEL: i = -276
# KERNEL: i = -277
# KERNEL: i = -278
# KERNEL: i = -279
# KERNEL: i = -280
# KERNEL: i = -281
# KERNEL: i = -282
# KERNEL: i = -283
# KERNEL: i = -284
# KERNEL: i = -285
# KERNEL: i = -286
# KERNEL: i = -287
# KERNEL: i = -288
# KERNEL: i = -289
# KERNEL: i = -290
# KERNEL: i = -291
# KERNEL: i = -292
# KERNEL: i = -293
# KERNEL: i = -294
# KERNEL: i = -295
# KERNEL: i = -296
# KERNEL: i = -297
# KERNEL: i = -298
# KERNEL: i = -299
# KERNEL: i = -300
# KERNEL: i = -301
# KERNEL: i = -302
# KERNEL: i = -303
# KERNEL: i = -304
# KERNEL: i = -305
# KERNEL: i = -306
# KERNEL: i = -307
# KERNEL: i = -308
# KERNEL: i = -309
# KERNEL: i = -310
# KERNEL: i = -311
# KERNEL: i = -312
# KERNEL: i = -313
# KERNEL: i = -314
# KERNEL: i = -315
# KERNEL: i = -316
# KERNEL: i = -317
# KERNEL: i = -318
# KERNEL: i = -319
# KERNEL: i = -320
# KERNEL: i = -321
# KERNEL: i = -322
# KERNEL: i = -323
# KERNEL: i = -324
# KERNEL: i = -325
# KERNEL: i = -326
# KERNEL: i = -327
# KERNEL: i = -328
# KERNEL: i = -329
# KERNEL: i = -330
# KERNEL: i = -331
# KERNEL: i = -332
# KERNEL: i = -333
# KERNEL: i = -334
# KERNEL: i = -335
# KERNEL: i = -336
# KERNEL: i = -337
# KERNEL: i = -338
# KERNEL: i = -339
# KERNEL: i = -340
# KERNEL: i = -341
# KERNEL: i = -342
# KERNEL: i = -343
# KERNEL: i = -344
# KERNEL: i = -345
# KERNEL: i = -346
# KERNEL: i = -347
# KERNEL: i = -348
# KERNEL: i = -349
# KERNEL: i = -350
# KERNEL: i = -351
# KERNEL: i = -352
# KERNEL: i = -353
# KERNEL: i = -354
# KERNEL: i = -355
# KERNEL: i = -356
# KERNEL: i = -357
# KERNEL: i = -358
# KERNEL: i = -359
# KERNEL: i = -360
# KERNEL: i = -361
# KERNEL: i = -362
# KERNEL: i = -363
# KERNEL: i = -364
# KERNEL: i = -365
# KERNEL: i = -366
# KERNEL: i = -367
# KERNEL: i = -368
# KERNEL: i = -369
# KERNEL: i = -370
# KERNEL: i = -371
# KERNEL: i = -372
# KERNEL: i = -373
# KERNEL: i = -374
# KERNEL: i = -375
# KERNEL: i = -376
# KERNEL: i = -377
# KERNEL: i = -378
# KERNEL: i = -379
# KERNEL: i = -380
# KERNEL: i = -381
# KERNEL: i = -382
# KERNEL: i = -383
# KERNEL: i = -384
# KERNEL: i = -385
# KERNEL: i = -386
# KERNEL: i = -387
# KERNEL: i = -388
# KERNEL: i = -389
# KERNEL: i = -390
# KERNEL: i = -391
# KERNEL: i = -392
# KERNEL: i = -393
# KERNEL: i = -394
# KERNEL: i = -395
# KERNEL: i = -396
# KERNEL: i = -397
# KERNEL: i = -398
# KERNEL: i = -399
# KERNEL: i = -400
# KERNEL: i = -401
# KERNEL: i = -402
# KERNEL: i = -403
# KERNEL: i = -404
# KERNEL: i = -405
# KERNEL: i = -406
# KERNEL: i = -407
# KERNEL: i = -408
# KERNEL: i = -409
# KERNEL: i = -410
# KERNEL: i = -411
# KERNEL: i = -412
# KERNEL: i = -413
# KERNEL: i = -414
# KERNEL: i = -415
# KERNEL: i = -416
# KERNEL: i = -417
# KERNEL: i = -418
# KERNEL: i = -419
# KERNEL: i = -420
# KERNEL: i = -421
# KERNEL: i = -422
# KERNEL: i = -423
# KERNEL: i = -424
# KERNEL: i = -425
# KERNEL: i = -426
# KERNEL: i = -427
# KERNEL: i = -428
# KERNEL: i = -429
# KERNEL: i = -430
# KERNEL: i = -431
# KERNEL: i = -432
# KERNEL: i = -433
# KERNEL: i = -434
# KERNEL: i = -435
# KERNEL: i = -436
# KERNEL: i = -437
# KERNEL: i = -438
# KERNEL: i = -439
# KERNEL: i = -440
# KERNEL: i = -441
# KERNEL: i = -442
# KERNEL: i = -443
# KERNEL: i = -444
# KERNEL: i = -445
# KERNEL: i = -446
# KERNEL: i = -447
# KERNEL: i = -448
# KERNEL: i = -449
# KERNEL: i = -450
# KERNEL: i = -451
# KERNEL: i = -452
# KERNEL: i = -453
# KERNEL: i = -454
# KERNEL: i = -455
# KERNEL: i = -456
# KERNEL: i = -457
# KERNEL: i = -458
# KERNEL: i = -459
# KERNEL: i = -460
# KERNEL: i = -461
# KERNEL: i = -462
# KERNEL: i = -463
# KERNEL: i = -464
# KERNEL: i = -465
# KERNEL: i = -466
# KERNEL: i = -467
# KERNEL: i = -468
# KERNEL: i = -469
# KERNEL: i = -470
# KERNEL: i = -471
# KERNEL: i = -472
# KERNEL: i = -473
# KERNEL: i = -474
# KERNEL: i = -475
# KERNEL: i = -476
# KERNEL: i = -477
# KERNEL: i = -478
# KERNEL: i = -479
# KERNEL: i = -480
# KERNEL: i = -481
# KERNEL: i = -482
# KERNEL: i = -483
# KERNEL: i = -484
# KERNEL: i = -485
# KERNEL: i = -486
# KERNEL: i = -487
# KERNEL: i = -488
# KERNEL: i = -489
# KERNEL: i = -490
# KERNEL: i = -491
# KERNEL: i = -492
# KERNEL: i = -493
# KERNEL: i = -494
# KERNEL: i = -495
# KERNEL: i = -496
# KERNEL: i = -497
# KERNEL: i = -498
# KERNEL: i = -499
# KERNEL: i = -500
# KERNEL: i = -501
# KERNEL: i = -502
# KERNEL: i = -503
# KERNEL: i = -504
# KERNEL: i = -505
# KERNEL: i = -506
# KERNEL: i = -507
# KERNEL: i = -508
# KERNEL: i = -509
# KERNEL: i = -510
# KERNEL: i = -511
# KERNEL: i = -512
# KERNEL: i = -513
# KERNEL: i = -514
# KERNEL: i = -515
# KERNEL: i = -516
# KERNEL: i = -517
# KERNEL: i = -518
# KERNEL: i = -519
# KERNEL: i = -520
# KERNEL: i = -521
# KERNEL: i = -522
# KERNEL: i = -523
# KERNEL: i = -524
# KERNEL: i = -525
# KERNEL: i = -526
# KERNEL: i = -527
# KERNEL: i = -528
# KERNEL: i = -529
# KERNEL: i = -530
# KERNEL: i = -531
# KERNEL: i = -532
# KERNEL: i = -533
# KERNEL: i = -534
# KERNEL: i = -535
# KERNEL: i = -536
# KERNEL: i = -537
# KERNEL: i = -538
# KERNEL: i = -539
# KERNEL: i = -540
# KERNEL: i = -541
# KERNEL: i = -542
# KERNEL: i = -543
# KERNEL: i = -544
# KERNEL: i = -545
# KERNEL: i = -546
# KERNEL: i = -547
# KERNEL: i = -548
# KERNEL: i = -549
# KERNEL: i = -550
# KERNEL: i = -551
# KERNEL: i = -552
# KERNEL: i = -553
# KERNEL: i = -554
# KERNEL: i = -555
# KERNEL: i = -556
# KERNEL: i = -557
# KERNEL: i = -558
# KERNEL: i = -559
# KERNEL: i = -560
# KERNEL: i = -561
# KERNEL: i = -562
# KERNEL: i = -563
# KERNEL: i = -564
# KERNEL: i = -565
# KERNEL: i = -566
# KERNEL: i = -567
# KERNEL: i = -568
# KERNEL: i = -569
# KERNEL: i = -570
# KERNEL: i = -571
# KERNEL: i = -572
# KERNEL: i = -573
# KERNEL: i = -574
# KERNEL: i = -575
# KERNEL: i = -576
# KERNEL: i = -577
# KERNEL: i = -578
# KERNEL: i = -579
# KERNEL: i = -580
# KERNEL: i = -581
# KERNEL: i = -582
# KERNEL: i = -583
# KERNEL: i = -584
# KERNEL: i = -585
# KERNEL: i = -586
# KERNEL: i = -587
# KERNEL: i = -588
# KERNEL: i = -589
goes to infinity.......
