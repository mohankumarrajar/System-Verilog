module forever_ex;
    initial begin
        forever begin
          $display("get the solution");
            #10;
          break;
          $display("
        end
    end
  initial begin
    $dumpfile("fuif.vcd");
    $dumpvars();
  end
  
endmodule


output :

                   get the solution
