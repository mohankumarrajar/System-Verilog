module ex4;
  string names[3] = '{"Mohankumar", "Divya", "Priya"};
  initial $display("Second name = %s", names[1]);
endmodule

output : Second name = Divya
