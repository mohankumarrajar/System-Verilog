module for_loop;
  
  initial begin
    
    for (int i = 0; i < 5;i ++)begin
      $display("putting the values the positve",i);
      
    end
  end
endmodule

output :

putting the values the positve          0
putting the values the positve          1
putting the values the positve          2
putting the values the positve          3
putting the values the positve          4
