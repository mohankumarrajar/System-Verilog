module ex1;
  logic [3:0] a;
  initial begin
    a = 4'b1010;
    $display("a = %b", a);
  end
endmodule
output : a = 1010
