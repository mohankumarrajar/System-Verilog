module m9;
  initial begin
    $display("Hello");
    repeat (3);
    
  end
endmodule

output :

# KERNEL: Hello
# KERNEL: Simulation has finished.
