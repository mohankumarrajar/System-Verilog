module m9;
  initial begin
    repeat (3) $display("Hello");
  end
endmodule


output :

# KERNEL: Hello
# KERNEL: Hello
# KERNEL: Hello
# KERNEL: Simulation has finished.
