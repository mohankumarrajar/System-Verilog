module tb;
	initial begin
		repeat (5) begin
			$display ("Repeat this statement");
		end
	end
endmodule

output : 
# KERNEL: Repeat this statement
# KERNEL: Repeat this statement
# KERNEL: Repeat this statement
# KERNEL: Repeat this statement
# KERNEL: Repeat this statement
# KERNEL: Simulation has finished
