module m1;
  int a;
  initial begin
    a = 1010;
    $display("a = %0d", a);
  end
endmodule

output :

# KERNEL: a = 1010
# KERNEL: Simulation has finished. 
